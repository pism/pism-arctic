netcdf pism_overrides {
    variables:
    byte pism_overrides;

    pism_overrides:grid.allow_extrapolation = "yes";

    pism_overrides:energy.minimum_allowed_temperature = 0.0;

    pism_overrides:stress_balance.sia.max_diffusivity = 100000.0;

    pism_overrides:surface.pdd.air_temp_all_precip_as_snow = 272.15;

    pism_overrides:surface.pdd.air_temp_all_precip_as_rain = 274.15;

    pism_overrides:surface.pdd.refreeze = 0.47;

    pism_overrides:surface.pdd.refreeze_ice_melt = "no";

    pism_overrides:run_info.institution = "University of Alaska Fairbanks";
    pism_overrides:run_info.institution_doc = "Institution name. This string is written to output files as the 'institution' global attribute.";

    pism_overrides:output.backup_interval = 5.0;
    pism_overrides:output.backup_interval_doc = "hours; wall-clock time between automatic backups";
    
    pism_overrides:surface.force_to_thickness.alpha = 0.1;
    pism_overrides:surface.force_to_thickness.alpha_doc = "yr-1; exponential coefficient in force-to-thickness mechanism";

    pism_overrides:surface.force_to_thickness.ice_free_alpha_factor = 5.0;
    pism_overrides:surface.force_to_thickness.ice_free_alpha_factor_doc = "; force_to_thickness_alpha is multiplied by this factor in areas that are ice-free according to the target ice thickness and force_to_thickness_ice_free_thickness_threshold";

    pism_overrides:ocean.sub_shelf_heat_flux_into_ice = 50.0;
    pism_overrides:ocean.sub_shelf_heat_flux_into_ice_doc = "W m-2; = J m-2 s-1; naively chosen default value for heat from ocean; see comments in @ref pism::POConstant::shelf_base_mass_flux().";

    pism_overrides:geometry.ice_free_thickness_standard = 10.0;

    pism_overrides:stress_balance.sia.bed_smoother.range = 5.0e2;

}
